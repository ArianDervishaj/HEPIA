--==============================================================================
--== Logisim goes FPGA automatic generated VHDL code                          ==
--==                                                                          ==
--==                                                                          ==
--== Project   : Add1bit                                                      ==
--== Component : Add1bit                                                      ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY Add1bit IS
   PORT ( A                         : IN  std_logic;
          B                         : IN  std_logic;
          C_in                      : IN  std_logic;
          C_out                     : OUT std_logic;
          D                         : OUT std_logic);
END Add1bit;

