--==============================================================================
--== Logisim goes FPGA automatic generated VHDL code                          ==
--==                                                                          ==
--==                                                                          ==
--== Project   : Add1bit                                                      ==
--== Component : LogisimToplevelShell                                         ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY LogisimToplevelShell IS
   PORT ( FPGA_INPUT_PIN_0          : IN  std_logic;
          FPGA_INPUT_PIN_1          : IN  std_logic;
          FPGA_INPUT_PIN_10         : IN  std_logic;
          FPGA_INPUT_PIN_11         : IN  std_logic;
          FPGA_INPUT_PIN_12         : IN  std_logic;
          FPGA_INPUT_PIN_13         : IN  std_logic;
          FPGA_INPUT_PIN_14         : IN  std_logic;
          FPGA_INPUT_PIN_15         : IN  std_logic;
          FPGA_INPUT_PIN_16         : IN  std_logic;
          FPGA_INPUT_PIN_2          : IN  std_logic;
          FPGA_INPUT_PIN_3          : IN  std_logic;
          FPGA_INPUT_PIN_4          : IN  std_logic;
          FPGA_INPUT_PIN_5          : IN  std_logic;
          FPGA_INPUT_PIN_6          : IN  std_logic;
          FPGA_INPUT_PIN_7          : IN  std_logic;
          FPGA_INPUT_PIN_8          : IN  std_logic;
          FPGA_INPUT_PIN_9          : IN  std_logic;
          FPGA_OUTPUT_PIN_0         : OUT std_logic;
          FPGA_OUTPUT_PIN_1         : OUT std_logic;
          FPGA_OUTPUT_PIN_2         : OUT std_logic;
          FPGA_OUTPUT_PIN_3         : OUT std_logic;
          FPGA_OUTPUT_PIN_4         : OUT std_logic;
          FPGA_OUTPUT_PIN_5         : OUT std_logic;
          FPGA_OUTPUT_PIN_6         : OUT std_logic;
          FPGA_OUTPUT_PIN_7         : OUT std_logic;
          FPGA_OUTPUT_PIN_8         : OUT std_logic);
END LogisimToplevelShell;

